// DEFINES
`define BITS 2         // Bit width of the operands

module 	bm_dag1_log(clock, 
		a_in, 
		b_in, 
		out);

// SIGNAL DECLARATIONS
input	clock;

input [`BITS-1:0] a_in;
input [`BITS-1:0] b_in;

output [`BITS-1:0] out;

wire [`BITS-1:0]    out;
wire [`BITS-1:0]    temp1;
wire [`BITS-1:0]    temp2;
wire [`BITS-1:0]    temp3;

// ASSIGN STATEMENTS
assign out = temp1 | temp2 | temp3;
assign temp1 = a_in & b_in;
assign temp2 = a_in ^ b_in;
assign temp3 = b_in ^ b_in;

endmodule
